`timescale 1ns/1ns

module InstructionMemory(
    input [31:0]address,
    output [31:0]instruction
); 
    reg [31:0] instructions [127:0];
	initial begin 
		instructions[0] = 32'b1110_00_1_1101_0_0000_0000_000000010100;
        instructions[1] = 32'b1110_00_1_1101_0_0000_0001_101000000001;
        instructions[2] = 32'b1110_00_1_1101_0_0000_0010_000100000011;
        instructions[3] = 32'b1110_00_0_0100_1_0010_0011_000000000010;
        instructions[4] = 32'b1110_00_0_0101_0_0000_0100_000000000000;
        instructions[5] = 32'b1110_00_0_0010_0_0100_0101_000100000100;
        instructions[6] = 32'b1110_00_0_0110_0_0000_0110_000010100000;
        instructions[7] = 32'b1110_00_0_1100_0_0101_0111_000101000010;
        instructions[8] = 32'b1110_00_0_0000_0_0111_1000_000000000011;
        instructions[9] = 32'b1110_00_0_1111_0_0000_1001_000000000110;
        instructions[10] = 32'b1110_00_0_0001_0_0100_1010_000000000101;
        instructions[11] = 32'b1110_00_0_1010_1_1000_0000_000000000110;
        instructions[12] = 32'b0001_00_0_0100_0_0001_0001_000000000001;
        instructions[13] = 32'b1110_00_0_1000_1_1001_0000_000000001000;
        instructions[14] = 32'b0000_00_0_0100_0_0010_0010_000000000010;
        instructions[15] = 32'b1110_00_1_1101_0_0000_0000_101100000001;
        instructions[16] = 32'b1110_01_0_0100_0_0000_0001_000000000000;
        instructions[17] = 32'b1110_01_0_0100_1_0000_1011_000000000000;
        instructions[18] = 32'b1110_01_0_0100_0_0000_0010_000000000100;
        instructions[19] = 32'b1110_01_0_0100_0_0000_0011_000000001000;
        instructions[20] = 32'b1110_01_0_0100_0_0000_0100_000000001101;
        instructions[21] = 32'b1110_01_0_0100_0_0000_0101_000000010000;
        instructions[22] = 32'b1110_01_0_0100_0_0000_0110_000000010100;
        instructions[23] = 32'b1110_01_0_0100_1_0000_1010_000000000100;
        instructions[24] = 32'b1110_01_0_0100_0_0000_0111_000000011000;
        instructions[25] = 32'b1110_00_1_1101_0_0000_0001_000000000100;
        instructions[26] = 32'b1110_00_1_1101_0_0000_0010_000000000000;
        instructions[27] = 32'b1110_00_1_1101_0_0000_0011_000000000000;
        instructions[28] = 32'b1110_00_0_0100_0_0000_0100_000100000011;
        instructions[29] = 32'b1110_01_0_0100_1_0100_0101_000000000000;
        instructions[30] = 32'b1110_01_0_0100_1_0100_0110_000000000100;
        instructions[31] = 32'b1110_00_0_1010_1_0101_0000_000000000110;
        instructions[32] = 32'b1100_01_0_0100_0_0100_0110_000000000000;
        instructions[33] = 32'b1100_01_0_0100_0_0100_0101_000000000100;
        instructions[34] = 32'b1110_00_1_0100_0_0011_0011_000000000001;
        instructions[35] = 32'b1110_00_1_1010_1_0011_0000_000000000011;
        instructions[36] = 32'b1011_10_1_0_111111111111111111110111;
        instructions[37] = 32'b1110_00_1_0100_0_0010_0010_000000000001;
        instructions[38] = 32'b1110_00_0_1010_1_0010_0000_000000000001;
        instructions[39] = 32'b1011_10_1_0_111111111111111111110011;
        instructions[40] = 32'b1110_01_0_0100_1_0000_0001_000000000000;
        instructions[41] = 32'b1110_01_0_0100_1_0000_0010_000000000100;
        instructions[42] = 32'b1110_01_0_0100_1_0000_0011_000000001000;
        instructions[43] = 32'b1110_01_0_0100_1_0000_0100_000000001100;
        instructions[44] = 32'b1110_01_0_0100_1_0000_0101_000000010000;
        instructions[45] = 32'b1110_01_0_0100_1_0000_0110_000000010100;
        instructions[46] = 32'b1110_10_1_0_111111111111111111111111;
	end
	assign instruction = instructions[address/4];
endmodule